library verilog;
use verilog.vl_types.all;
entity Integrador_vlg_vec_tst is
end Integrador_vlg_vec_tst;
